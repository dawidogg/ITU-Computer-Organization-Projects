module control_unit_tb;

  reg clk;
  control_unit uut(clk);
  
  
  initial begin
    clk = 0;
  end
endmodule